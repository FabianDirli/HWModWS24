library ieee;
use ieee.std_logic_1164.all;
use work.sram_ctrl_pkg.all;
package test_sequence_pkg is
	constant TEST_SEQUENCE : sequence_t := (x"1313",x"0CCE",x"8CD0",x"7D62",x"7248",x"4771",x"347A",x"2C83",x"D806",x"1045",x"0F41",x"2FF8",x"6FF1",x"771F",x"0D96",x"65CE",x"6574",x"765F",x"76C6",x"86C1",x"7202",x"264D",x"26FF",x"56E6",x"265D",x"72C2",x"8205",x"762D",x"7752",x"7740",x"8201",x"274D",x"8681",x"7615",x"7746",x"8270",x"273D",x"8201",x"76EC",x"26FD",x"674F",x"7202",x"261D",x"76C5",x"66CE",x"73AF",x"7201",x"7492",x"76EF",x"220D",x"76D6",x"779B",x"220D",x"5721",x"5651",x"56D0",x"461E",x"269E",x"26EF",x"273D",x"8201",x"779C",x"26FD",x"775C",x"8202",x"773F",x"268D",x"761A",x"66CE",x"76C6",x"7209",x"266D",x"8691",x"76EC",x"264D",x"7204",x"674E",x"7686",x"761B",x"274D",x"620E",x"261D",x"620F",x"772C",x"76FB",x"86D2",x"8610",x"26ED",x"720D",x"765C",x"76D6",x"770B",x"8651",x"372B",x"26FD",x"572A",x"620E",x"7688",x"7612",x"273D",x"8200",x"8682",x"769F",x"7642",x"264D",x"8651",x"76EC",x"220D",x"677E",x"7689",x"8610",x"774C",x"220D",x"679E",x"86F1",x"8751",x"620E",x"7730",x"7655",x"265D",x"86B6",x"720C",x"86F2",x"76EF",x"220D",x"7610",x"720C",x"7641",x"7612",x"279D",x"720D",x"76FF",x"766C",x"7201",x"86D2",x"7690",x"7736",x"766B",x"76F4",x"272D",x"8741",x"7755",x"76E6",x"8650",x"32EB",x"D6CB",x"70DD",x"E5FE",x"8E6F",x"0353",x"51BE",x"D860",x"AE35",x"8E45",x"4F9B",x"6E3D",x"AC56",x"3454",x"2F7C",x"C285",x"3184");
end package;
